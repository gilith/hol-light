/*----------------------------------------------------------------------------+
| module montgomery91 satisfies the following property:                       |
|                                                                             |
| !x y t.                                                                     |
|     (!i. i <= 12 ==> (signal ld (t + i) <=> i = 0)) /\                      |
|     bits_to_num (bsignal xs[0:6] t) + 2 * bits_to_num (bsignal xc[0:6] t) = |
|     x /\                                                                    |
|     (!i. 2 <= i /\ i <= 10                                                  |
|          ==> bits_to_num (bsignal ys[0:6] (t + i)) +                        |
|              2 * bits_to_num (bsignal yc[0:6] (t + i)) =                    |
|              y)                                                             |
|     ==> bits_to_num (bsignal zs[0:7] (t + 15)) +                            |
|         2 * bits_to_num (bsignal zc[0:7] (t + 15)) =                        |
|         montgomery_reduce 91 (2 EXP 9) 45 (x * y)                           |
+----------------------------------------------------------------------------*/

module montgomery91(clk,ld,xs,xc,ys,yc,zs,zc);
  input clk;
  input ld;
  input [0:6] xs;
  input [0:6] xc;
  input [0:6] ys;
  input [0:6] yc;

  output [0:7] zs;
  output [0:7] zc;

  reg r0;
  reg r1;
  reg r2;
  reg r3;
  reg r4;
  reg r5;
  reg r6;
  reg r7;
  reg r8;
  reg r9;
  reg r10;
  reg r11;
  reg r12;
  reg r13;
  reg r14;
  reg r15;
  reg r16;
  reg r17;
  reg r18;
  reg r19;
  reg r20;
  reg r21;
  reg r22;
  reg r23;
  reg r24;
  reg r25;
  reg r26;
  reg r27;
  reg r28;
  reg r29;
  reg r30;
  reg r31;
  reg r32;
  reg r33;
  reg r34;
  reg r35;
  reg r36;
  reg r37;
  reg r38;
  reg r39;
  reg r40;
  reg r41;
  reg r42;
  reg r43;
  reg r44;
  reg r45;
  reg r46;
  reg r47;
  reg r48;
  reg r49;
  reg r50;
  reg r51;
  reg r52;
  reg r53;
  reg r54;
  reg r55;
  reg r56;
  reg r57;
  reg r58;
  reg r59;
  reg r60;
  reg r61;
  reg r62;
  reg r63;
  reg r64;
  reg r65;
  reg r66;
  reg r67;
  reg r68;
  reg r69;

  wire w0;
  wire w1;
  wire w2;
  wire w3;
  wire w4;
  wire w5;
  wire w6;
  wire w7;
  wire w8;
  wire w9;
  wire w10;
  wire w11;
  wire w12;
  wire w13;
  wire w14;
  wire w15;
  wire w16;
  wire w17;
  wire w18;
  wire w19;
  wire w20;
  wire w21;
  wire w22;
  wire w23;
  wire w24;
  wire w25;
  wire w26;
  wire w27;
  wire w28;
  wire w29;
  wire w30;
  wire w31;
  wire w32;
  wire w33;
  wire w34;
  wire w35;
  wire w36;
  wire w37;
  wire w38;
  wire w39;
  wire w40;
  wire w41;
  wire w42;
  wire w43;
  wire w44;
  wire w45;
  wire w46;
  wire w47;
  wire w48;
  wire w49;
  wire w50;
  wire w51;
  wire w52;
  wire w53;
  wire w54;
  wire w55;
  wire w56;
  wire w57;
  wire w58;
  wire w59;
  wire w60;
  wire w61;
  wire w62;
  wire w63;
  wire w64;
  wire w65;
  wire w66;
  wire w67;
  wire w68;
  wire w69;
  wire w70;
  wire w71;
  wire w72;
  wire w73;
  wire w74;
  wire w75;
  wire w76;
  wire w77;
  wire w78;
  wire w79;
  wire w80;
  wire w81;
  wire w82;
  wire w83;
  wire w84;
  wire w85;
  wire w86;
  wire w87;
  wire w88;
  wire w89;
  wire w90;
  wire w91;
  wire w92;
  wire w93;
  wire w94;
  wire w95;
  wire w96;
  wire w97;
  wire w98;
  wire w99;
  wire w100;
  wire w101;
  wire w102;
  wire w103;
  wire w104;
  wire w105;
  wire w106;
  wire w107;
  wire w108;
  wire w109;
  wire w110;
  wire w111;
  wire w112;
  wire w113;
  wire w114;
  wire w115;
  wire w116;
  wire w117;
  wire w118;
  wire w119;
  wire w120;
  wire w121;
  wire w122;
  wire w123;
  wire w124;
  wire w125;
  wire w126;
  wire w127;
  wire w128;
  wire w129;
  wire w130;
  wire w131;
  wire w132;
  wire w133;
  wire w134;
  wire w135;
  wire w136;
  wire w137;
  wire w138;
  wire w139;
  wire w140;
  wire w141;
  wire w142;
  wire w143;
  wire w144;
  wire w145;
  wire w146;
  wire w147;
  wire w148;
  wire w149;
  wire w150;
  wire w151;
  wire w152;
  wire w153;
  wire w154;
  wire w155;
  wire w156;
  wire w157;
  wire w158;
  wire w159;
  wire w160;
  wire w161;
  wire w162;
  wire w163;
  wire w164;
  wire w165;
  wire w166;
  wire w167;
  wire w168;
  wire w169;
  wire w170;
  wire w171;
  wire w172;
  wire w173;
  wire w174;
  wire w175;
  wire w176;
  wire w177;
  wire w178;
  wire w179;
  wire w180;
  wire w181;
  wire w182;
  wire w183;
  wire w184;
  wire w185;
  wire w186;
  wire w187;
  wire w188;
  wire w189;
  wire w190;
  wire w191;
  wire w192;
  wire w193;
  wire w194;
  wire w195;
  wire w196;
  wire w197;
  wire w198;
  wire w199;
  wire w200;
  wire w201;
  wire w202;
  wire w203;
  wire w204;
  wire w205;
  wire w206;
  wire w207;
  wire w208;
  wire w209;
  wire w210;
  wire w211;
  wire w212;
  wire w213;
  wire w214;
  wire w215;
  wire w216;
  wire w217;
  wire w218;
  wire w219;
  wire w220;
  wire w221;
  wire w222;
  wire w223;
  wire w224;
  wire w225;
  wire w226;
  wire w227;
  wire w228;
  wire w229;
  wire w230;
  wire w231;
  wire w232;
  wire w233;
  wire w234;
  wire w235;
  wire w236;
  wire w237;
  wire w238;
  wire w239;
  wire w240;
  wire w241;
  wire w242;
  wire w243;
  wire w244;
  wire w245;
  wire w246;
  wire w247;
  wire w248;
  wire w249;
  wire w250;
  wire w251;
  wire w252;
  wire w253;
  wire w254;
  wire w255;
  wire w256;
  wire w257;
  wire w258;
  wire w259;
  wire w260;
  wire w261;
  wire w262;
  wire w263;
  wire w264;
  wire w265;
  wire w266;
  wire w267;
  wire w268;
  wire w269;
  wire w270;
  wire w271;
  wire w272;
  wire w273;
  wire w274;
  wire w275;
  wire w276;
  wire w277;
  wire w278;
  wire w279;
  wire w280;
  wire w281;
  wire w282;
  wire w283;
  wire w284;
  wire w285;
  wire w286;
  wire w287;
  wire w288;
  wire w289;
  wire w290;
  wire w291;
  wire w292;
  wire w293;
  wire w294;
  wire w295;
  wire w296;
  wire w297;
  wire w298;
  wire w299;
  wire w300;
  wire w301;
  wire w302;
  wire w303;
  wire w304;
  wire w305;
  wire w306;
  wire w307;
  wire w308;
  wire w309;
  wire w310;
  wire w311;
  wire w312;
  wire w313;
  wire w314;
  wire w315;
  wire w316;
  wire w317;
  wire w318;
  wire w319;
  wire w320;
  wire w321;
  wire w322;
  wire w323;
  wire w324;
  wire w325;
  wire w326;
  wire w327;
  wire w328;
  wire w329;
  wire w330;
  wire w331;
  wire w332;
  wire w333;
  wire w334;
  wire w335;
  wire w336;
  wire w337;
  wire w338;
  wire w339;

  assign w0 = ld ? xs[6] : r0;
  assign w1 = ld ? xs[5] : w2;
  assign w2 = r12 ^ r11;
  assign w3 = ld ? xs[4] : w4;
  assign w4 = r14 ^ r13;
  assign w5 = ld ? xs[3] : w6;
  assign w6 = r16 ^ r15;
  assign w7 = ld ? xs[2] : w8;
  assign w8 = r18 ^ r17;
  assign w9 = ld ? xs[1] : w10;
  assign w10 = r20 ^ r19;
  assign w11 = ld ? xs[0] : w12;
  assign w12 = r22 ^ r21;
  assign w13 = ld ? xc[5] : w14;
  assign w14 = r12 & r11;
  assign w15 = ld ? xc[4] : w16;
  assign w16 = r14 & r13;
  assign w17 = ld ? xc[3] : w18;
  assign w18 = r16 & r15;
  assign w19 = ld ? xc[2] : w20;
  assign w20 = r18 & r17;
  assign w21 = ld ? xc[1] : w22;
  assign w22 = r20 & r19;
  assign w23 = ld ? xc[0] : w24;
  assign w24 = r22 & r21;
  assign w25 = w27 ^ w26;
  assign w26 = w219 | w218;
  assign w27 = w73 ^ w43;
  assign w28 = w30 ^ w29;
  assign w29 = w221 | w220;
  assign w30 = w74 ^ w46;
  assign w31 = w33 ^ w32;
  assign w32 = w223 | w222;
  assign w33 = w75 ^ w49;
  assign w34 = w36 ^ w35;
  assign w35 = w225 | w224;
  assign w36 = w76 ^ w52;
  assign w37 = w39 ^ w38;
  assign w38 = w227 | w226;
  assign w39 = w77 ^ w55;
  assign w40 = w42 ^ w41;
  assign w41 = w93 & w92;
  assign w42 = w78 ^ w58;
  assign w43 = w45 ^ w44;
  assign w44 = r45 & ys[6];
  assign w45 = w80 ^ w79;
  assign w46 = w48 ^ w47;
  assign w47 = r45 & ys[5];
  assign w48 = w82 ^ w81;
  assign w49 = w51 ^ w50;
  assign w50 = r45 & ys[4];
  assign w51 = w84 ^ w83;
  assign w52 = w54 ^ w53;
  assign w53 = r45 & ys[3];
  assign w54 = w86 ^ w85;
  assign w55 = w57 ^ w56;
  assign w56 = r45 & ys[2];
  assign w57 = w88 ^ w87;
  assign w58 = w60 ^ w59;
  assign w59 = r45 & ys[1];
  assign w60 = w90 ^ w89;
  assign w61 = w63 ^ w62;
  assign w62 = w217 | w216;
  assign w63 = w72 ^ w71;
  assign w64 = r2 ^ r1;
  assign w65 = r3 ^ w66;
  assign w66 = r6 ^ r5;
  assign w67 = r4 ^ w68;
  assign w68 = w69 ^ r25;
  assign w69 = r8 ^ r7;
  assign w70 = r10 ^ r9;
  assign w71 = w322 & r40;
  assign w72 = r45 & yc[6];
  assign w73 = r45 & yc[5];
  assign w74 = r45 & yc[4];
  assign w75 = r45 & yc[3];
  assign w76 = r45 & yc[2];
  assign w77 = r45 & yc[1];
  assign w78 = r45 & yc[0];
  assign w79 = w322 & r41;
  assign w80 = w322 & r43;
  assign w81 = w322 & r42;
  assign w82 = w322 & r44;
  assign w83 = w322 & r39;
  assign w84 = w322 & r38;
  assign w85 = w322 & r2;
  assign w86 = w322 & r1;
  assign w87 = w322 & r3;
  assign w88 = w322 & r6;
  assign w89 = w322 & r4;
  assign w90 = w322 & r8;
  assign w91 = w93 ^ w92;
  assign w92 = r45 & ys[0];
  assign w93 = w322 & r10;
  assign w94 = w96 ^ w95;
  assign w95 = w118 & w117;
  assign w96 = w116 ^ w115;
  assign w97 = w99 ^ w98;
  assign w98 = w247 | w246;
  assign w99 = w118 ^ w117;
  assign w100 = w101 ^ r23;
  assign w101 = w120 ^ w119;
  assign w102 = w104 ^ w103;
  assign w103 = w249 | w248;
  assign w104 = w122 ^ w121;
  assign w105 = w106 ^ r23;
  assign w106 = w124 ^ w123;
  assign w107 = w108 ^ r23;
  assign w108 = w126 ^ w125;
  assign w109 = w111 ^ w110;
  assign w110 = w130 & r23;
  assign w111 = w128 ^ w127;
  assign w112 = w114 ^ w113;
  assign w113 = w116 & w115;
  assign w114 = w327 & r46;
  assign w115 = w327 & r47;
  assign w116 = w327 & r54;
  assign w117 = w327 & r48;
  assign w118 = w327 & r55;
  assign w119 = w327 & r49;
  assign w120 = w327 & r56;
  assign w121 = w327 & r50;
  assign w122 = w327 & r57;
  assign w123 = w327 & r51;
  assign w124 = w327 & r58;
  assign w125 = w327 & r52;
  assign w126 = w327 & r59;
  assign w127 = w327 & r53;
  assign w128 = w327 & r60;
  assign w129 = w130 ^ r23;
  assign w130 = w327 & r61;
  assign w131 = w100 ^ w132;
  assign w132 = w122 & w121;
  assign w133 = w105 ^ w134;
  assign w134 = w251 | w250;
  assign w135 = w107 ^ w136;
  assign w136 = w128 & w127;
  assign w137 = w139 ^ w138;
  assign w138 = w259 | w258;
  assign w139 = w153 ^ w152;
  assign w140 = w141 ^ r24;
  assign w141 = w155 ^ w154;
  assign w142 = w143 ^ r24;
  assign w143 = w157 ^ w156;
  assign w144 = w146 ^ w145;
  assign w145 = w263 | w262;
  assign w146 = w159 ^ w158;
  assign w147 = w148 ^ r24;
  assign w148 = w161 ^ w160;
  assign w149 = w151 ^ w150;
  assign w150 = w153 & w152;
  assign w151 = r24 ^ w185;
  assign w152 = w334 & r25;
  assign w153 = w334 & r7;
  assign w154 = w334 & r26;
  assign w155 = w334 & r9;
  assign w156 = w334 & r27;
  assign w157 = w334 & r36;
  assign w158 = w334 & r28;
  assign w159 = w334 & r35;
  assign w160 = w334 & r29;
  assign w161 = w334 & r33;
  assign w162 = w163 ^ r24;
  assign w163 = w334 & r31;
  assign w164 = w140 ^ w165;
  assign w165 = w261 | w260;
  assign w166 = w142 ^ w167;
  assign w167 = w159 & w158;
  assign w168 = w147 ^ w169;
  assign w169 = w163 & r24;
  assign w170 = w70 ^ r26;
  assign w171 = w172 ^ r27;
  assign w172 = r37 ^ r36;
  assign w173 = w174 ^ r28;
  assign w174 = r23 ^ r35;
  assign w175 = w176 ^ r29;
  assign w176 = r34 ^ r33;
  assign w177 = w178 ^ r30;
  assign w178 = r32 ^ r31;
  assign w179 = w65 ^ w180;
  assign w180 = w276 | w275;
  assign w181 = w67 ^ w182;
  assign w182 = w278 | w277;
  assign w183 = w64 ^ w184;
  assign w184 = r6 & r5;
  assign w185 = w334 & r5;
  assign w186 = w188 | w187;
  assign w187 = w43 & w26;
  assign w188 = w205 | w204;
  assign w189 = w191 | w190;
  assign w190 = w46 & w29;
  assign w191 = w207 | w206;
  assign w192 = w194 | w193;
  assign w193 = w49 & w32;
  assign w194 = w209 | w208;
  assign w195 = w197 | w196;
  assign w196 = w52 & w35;
  assign w197 = w211 | w210;
  assign w198 = w200 | w199;
  assign w199 = w55 & w38;
  assign w200 = w213 | w212;
  assign w201 = w203 | w202;
  assign w202 = w58 & w41;
  assign w203 = w215 | w214;
  assign w204 = w73 & w26;
  assign w205 = w73 & w43;
  assign w206 = w74 & w29;
  assign w207 = w74 & w46;
  assign w208 = w75 & w32;
  assign w209 = w75 & w49;
  assign w210 = w76 & w35;
  assign w211 = w76 & w52;
  assign w212 = w77 & w38;
  assign w213 = w77 & w55;
  assign w214 = w78 & w41;
  assign w215 = w78 & w58;
  assign w216 = w79 & w44;
  assign w217 = w229 | w228;
  assign w218 = w81 & w47;
  assign w219 = w231 | w230;
  assign w220 = w83 & w50;
  assign w221 = w233 | w232;
  assign w222 = w85 & w53;
  assign w223 = w235 | w234;
  assign w224 = w87 & w56;
  assign w225 = w237 | w236;
  assign w226 = w89 & w59;
  assign w227 = w239 | w238;
  assign w228 = w80 & w44;
  assign w229 = w80 & w79;
  assign w230 = w82 & w47;
  assign w231 = w82 & w81;
  assign w232 = w84 & w50;
  assign w233 = w84 & w83;
  assign w234 = w86 & w53;
  assign w235 = w86 & w85;
  assign w236 = w88 & w56;
  assign w237 = w88 & w87;
  assign w238 = w90 & w59;
  assign w239 = w90 & w89;
  assign w240 = w242 | w241;
  assign w241 = w71 & w62;
  assign w242 = w244 | w243;
  assign w243 = w72 & w62;
  assign w244 = w72 & w71;
  assign w245 = r39 | r38;
  assign w246 = w119 & r23;
  assign w247 = w253 | w252;
  assign w248 = w123 & r23;
  assign w249 = w255 | w254;
  assign w250 = w125 & r23;
  assign w251 = w257 | w256;
  assign w252 = w120 & r23;
  assign w253 = w120 & w119;
  assign w254 = w124 & r23;
  assign w255 = w124 & w123;
  assign w256 = w126 & r23;
  assign w257 = w126 & w125;
  assign w258 = w154 & r24;
  assign w259 = w265 | w264;
  assign w260 = w156 & r24;
  assign w261 = w267 | w266;
  assign w262 = w160 & r24;
  assign w263 = w269 | w268;
  assign w264 = w155 & r24;
  assign w265 = w155 & w154;
  assign w266 = w157 & r24;
  assign w267 = w157 & w156;
  assign w268 = w161 & r24;
  assign w269 = w161 & w160;
  assign w270 = w272 | w271;
  assign w271 = w185 & w150;
  assign w272 = w274 | w273;
  assign w273 = r24 & w150;
  assign w274 = r24 & w185;
  assign w275 = r7 & r25;
  assign w276 = w292 | w291;
  assign w277 = r9 & r26;
  assign w278 = w294 | w293;
  assign w279 = w281 | w280;
  assign w280 = r36 & r27;
  assign w281 = w296 | w295;
  assign w282 = w284 | w283;
  assign w283 = r35 & r28;
  assign w284 = w298 | w297;
  assign w285 = w287 | w286;
  assign w286 = r33 & r29;
  assign w287 = w300 | w299;
  assign w288 = w290 | w289;
  assign w289 = r31 & r30;
  assign w290 = w302 | w301;
  assign w291 = r8 & r25;
  assign w292 = r8 & r7;
  assign w293 = r10 & r26;
  assign w294 = r10 & r9;
  assign w295 = r37 & r27;
  assign w296 = r37 & r36;
  assign w297 = r23 & r28;
  assign w298 = r23 & r35;
  assign w299 = r34 & r29;
  assign w300 = r34 & r33;
  assign w301 = r32 & r30;
  assign w302 = r32 & r31;
  assign w303 = w305 | w304;
  assign w304 = w66 & w180;
  assign w305 = w310 | w309;
  assign w306 = w308 | w307;
  assign w307 = w68 & w182;
  assign w308 = w312 | w311;
  assign w309 = r3 & w180;
  assign w310 = r3 & w66;
  assign w311 = r4 & w182;
  assign w312 = r4 & w68;
  assign w313 = w315 | w314;
  assign w314 = r1 & w184;
  assign w315 = w317 | w316;
  assign w316 = r2 & w184;
  assign w317 = r2 & r1;
  assign w318 = w245 | w313;
  assign w319 = w162 | w320;
  assign w320 = w334 & r30;
  assign w321 = ld & xc[6];
  assign w322 = ~r62;
  assign w323 = w96 & w95;
  assign w324 = w99 & w98;
  assign w325 = w104 & w103;
  assign w326 = w111 & w110;
  assign w327 = ~r63;
  assign w328 = w114 & w113;
  assign w329 = w100 & w132;
  assign w330 = w105 & w134;
  assign w331 = w107 & w136;
  assign w332 = w139 & w138;
  assign w333 = w146 & w145;
  assign w334 = ~r64;
  assign w335 = w140 & w165;
  assign w336 = w142 & w167;
  assign w337 = w147 & w169;
  assign w338 = ~r24;
  assign w339 = ~r23;
  assign zs[0] = w177;
  assign zs[1] = w175;
  assign zs[2] = w173;
  assign zs[3] = w171;
  assign zs[4] = w170;
  assign zs[5] = w181;
  assign zs[6] = w179;
  assign zs[7] = w183;
  assign zc[0] = w288;
  assign zc[1] = w285;
  assign zc[2] = w282;
  assign zc[3] = w279;
  assign zc[4] = 1'b0;
  assign zc[5] = w306;
  assign zc[6] = w303;
  assign zc[7] = w318;

  always @(posedge clk)
    begin
      r0 <= w321;
      r1 <= w31;
      r2 <= w195;
      r3 <= w198;
      r4 <= w201;
      r5 <= w270;
      r6 <= w34;
      r7 <= w149;
      r8 <= w37;
      r9 <= w137;
      r10 <= w40;
      r11 <= w13;
      r12 <= w0;
      r13 <= w15;
      r14 <= w1;
      r15 <= w17;
      r16 <= w3;
      r17 <= w19;
      r18 <= w5;
      r19 <= w21;
      r20 <= w7;
      r21 <= w23;
      r22 <= w9;
      r23 <= r37;
      r24 <= r69;
      r25 <= w332;
      r26 <= w335;
      r27 <= w336;
      r28 <= w333;
      r29 <= w337;
      r30 <= w319;
      r31 <= w168;
      r32 <= r34;
      r33 <= w144;
      r34 <= r23;
      r35 <= w166;
      r36 <= w164;
      r37 <= w91;
      r38 <= w28;
      r39 <= w192;
      r40 <= w240;
      r41 <= w186;
      r42 <= w189;
      r43 <= w61;
      r44 <= w25;
      r45 <= r67;
      r46 <= w328;
      r47 <= w323;
      r48 <= w324;
      r49 <= w329;
      r50 <= w325;
      r51 <= w330;
      r52 <= w331;
      r53 <= w326;
      r54 <= w112;
      r55 <= w94;
      r56 <= w97;
      r57 <= w131;
      r58 <= w102;
      r59 <= w133;
      r60 <= w135;
      r61 <= w109;
      r62 <= r65;
      r63 <= r66;
      r64 <= r68;
      r65 <= ld;
      r66 <= r62;
      r67 <= w11;
      r68 <= r63;
      r69 <= w129;
    end

endmodule // montgomery91
